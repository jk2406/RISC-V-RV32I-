// RV32I 5-Stage Pipelined CPU 

`timescale 1ns/1ps
module riscv_pipelined #(
    parameter XLEN = 32,
    parameter IMEM_WORDS = 1024,
    parameter DMEM_WORDS = 1024
)(
    input  logic              clk,
    input  logic              rst_p ,    // active high reset
    output logic dummy_out //Since this cpu doesn't have any output,to make code synthesizable a dummy output has been provided
);
    logic dummy_var=1'b1;//Dummy output always one
    assign dummy_out=dummy_var;
    
    
     logic [31:0] imem [0:IMEM_WORDS-1];
     logic [31:0] dmem [0:DMEM_WORDS-1];
     logic [31:0] imem_dout; // instruction memory output from IP BRAM block
     logic [31:0] dmem_dout; // data memory output from IP BRAM block

     logic [31:0] pc_addr;
    logic [31:0] dmem_addr;
    logic [31:0] pc;
    assign pc_addr   = pc[31:2];             // word-address for instruction memory
    logic [9:0] pc_addr_ip;
    logic [9:0] dmem_addr_ip;

    assign pc_addr_ip   = pc[11:2];             
    
    logic [31:0] ex_mem_wdata; //Declared ahead because it is used in BRAM(commented out)
    logic ex_mem_mem_we;
    logic [31:0] regs [0:31];
  
//-----------------------------------------------
//Following is the default IP block generated.This is autogenerated by vivado 
//  blk_mem_gen_0_wrapper u_imem ( 
//     // Port A: Instruction memory (read-only)
//     .clka(clk),
//     .ena(1'b1),
//     .wea(1'b0),           // no writes
//     .addra(pc_addr_ip),
//     .dina(32'b0),
//     .douta(imem_dout),

//     // Port B: Data memory (read/write)
//     .clkb(clk),
//     .enb(ex_mem_mem_we),   // enable write
//     .web(ex_mem_mem_we),
//     .addrb(dmem_addr_ip),
//     .dinb(ex_mem_wdata),
//     .doutb(dmem_dout)
// );

//FOllowing is the ILA(Integrated Logic Analyser) to tap pc(autogenerated by vivado)
//     ila_0 u_ila (
//     .clk(clk),            // connect the same clock as your CPU
//     .probe0(pc[31:0])      // 32-bit probe for your program counter
// //    .trig_out_ack(1'b1)
// );

    
 

   
    // --- Pipeline Register Definitions ---
    // IF/ID Register
    logic [31:0] if_id_instr;
    logic [31:0] if_id_pc;
    
    // ID/EX Register
    logic [31:0] id_ex_instr;
    logic [31:0] id_ex_pc;
    logic [31:0] id_ex_rdata1;
    logic [31:0] id_ex_rdata2;
    logic [31:0] id_ex_imm;
    logic [3:0]  id_ex_alu_op; // Expanded to handle all ALU ops
    logic id_ex_reg_we;
    logic id_ex_is_load, id_ex_is_store; 
    logic id_ex_is_branch, id_ex_is_jal, id_ex_is_jalr; 
    logic id_ex_is_rtype, id_ex_is_itype_alu;
    logic [4:0] id_ex_rs1, id_ex_rs2; 
    logic [4:0] id_ex_rd;
    
    // EX/MEM Register
    logic [31:0] ex_mem_pc_plus_4; 
    logic [31:0] ex_mem_alu_out;
    
    logic [4:0]  ex_mem_rd; 
    logic ex_mem_reg_we; 
    
    logic ex_mem_is_load;
    logic ex_mem_is_jal; 
    
    // MEM/WB Register
    logic [31:0] mem_wb_alu_out;
    logic [31:0] mem_wb_mem_rdata;
    logic [31:0] mem_wb_pc_plus_4;
    logic [4:0]  mem_wb_rd;
    logic mem_wb_reg_we; 
    logic mem_wb_is_load;
    logic mem_wb_is_jal;
    
    // --- Hazard Control Signals ---
    logic [1:0] forward_a; 
    logic [1:0] forward_b; 
    logic pc_stall;         // Data Hazard (Load-Use) Stall: Freezes PC/IF/ID
    logic id_ex_bubble;     // Data Hazard (Load-Use) Bubble: NOPs ID/EX
    logic ex_branch_taken;  // Control Hazard Resolution: Branch/Jump Taken
    logic [31:0] ex_branch_target; // Calculated branch/jump target address
    
    // --- ALU Operation Codes (4-bit) ---
    localparam ALU_ADD  = 4'h0;
    localparam ALU_SUB  = 4'h1;
    localparam ALU_SLL  = 4'h2;
    localparam ALU_SLT  = 4'h3;
    localparam ALU_SLTU = 4'h4;
    localparam ALU_XOR  = 4'h5;
    localparam ALU_SRL  = 4'h6;
    localparam ALU_SRA  = 4'h7;
    localparam ALU_OR   = 4'h8;
    localparam ALU_AND  = 4'h9;

    // =========================================================================
    // STAGE 1: INSTRUCTION FETCH (IF)
    // =========================================================================



    wire [31:0] instr_if = imem_dout;
    always_ff @(posedge clk or posedge rst_p) begin
        if (rst_p) pc <= 32'd0;
       
        else if (ex_branch_taken) begin
            pc <= ex_branch_target;
        end

        else if (pc_stall) begin
            pc <= pc; // PC holds its value(stalling)
        end
        // Default: PC increments by 4 (Predict Not Taken)
        else begin
            pc <= pc + 4;
        end
    end

    // IF/ID Register Update (Handles Control Hazard Flush and Data Hazard Stall)
    always_ff @(posedge clk or posedge rst_p) begin
        if (rst_p) begin
            if_id_instr <= 32'b0;
            if_id_pc    <= 32'b0;
        end 
        // FLUSH: If a branch/jump is taken, flush the IF/ID register to NOP.
        else if (ex_branch_taken) begin
            if_id_instr <= 32'b0; 
            if_id_pc    <= 32'b0;
        end 
        // STALL: If stalling, IF/ID holds its value.
        else if (pc_stall) begin
            if_id_instr <= if_id_instr; 
            if_id_pc    <= if_id_pc;    
        end
        // NORMAL: Pass instruction from IF to ID
        else begin
            if_id_instr <= instr_if;
            if_id_pc    <= pc;
        end
    end


    // =========================================================================
    // STAGE 2: INSTRUCTION DECODE / REGISTER FETCH (ID)
    // =========================================================================
    
  
    wire [6:0]  id_opcode = if_id_instr[6:0];
    wire [4:0]  id_rd     = if_id_instr[11:7];
    wire [2:0]  id_funct3 = if_id_instr[14:12];
    wire [4:0]  id_rs1    = if_id_instr[19:15];
    wire [4:0]  id_rs2    = if_id_instr[24:20];
    wire [6:0]  id_funct7 = if_id_instr[31:25];
    

    wire [31:0] id_rdata1 = (id_rs1 == 0) ? 32'b0 : regs[id_rs1];
    wire [31:0] id_rdata2 = (id_rs2 == 0) ? 32'b0 : regs[id_rs2];

    // Immediate Generation 
    wire [31:0] id_imm_i = {{20{if_id_instr[31]}}, if_id_instr[31:20]};
    wire [31:0] id_imm_s = {{20{if_id_instr[31]}}, if_id_instr[31:25], if_id_instr[11:7]};
    wire [31:0] id_imm_u_shifted = {if_id_instr[31:12], 12'b0};
    wire [31:0] id_imm_b; 
    wire [31:0] id_imm_j;

    // Branch Immediate (B-type)
   
    assign id_imm_b = {{19{if_id_instr[31]}}, if_id_instr[31:20],1'b0};//Last bit must be zero(even)
    
    // JAL Immediate (J-type)
  
    assign id_imm_j = {{12{if_id_instr[31]}}, if_id_instr[31:12]};
    
    // Control Unit- DECODING ALL ALU OPS
    logic id_reg_we;
    logic id_is_load, id_is_store, id_is_branch, id_is_jal, id_is_jalr;
    logic id_is_rtype, id_is_itype_alu;
    logic [3:0] id_alu_op;
    
    always_comb begin
        id_reg_we = 1'b0;
        id_is_load = 1'b0; id_is_store = 1'b0; id_is_branch = 1'b0; id_is_jal = 1'b0; id_is_jalr = 1'b0;
        id_is_rtype = 1'b0; id_is_itype_alu = 1'b0;
        id_alu_op = ALU_ADD; //For safety,defaulted to ADD

        unique case (id_opcode)
            7'b0110011: begin // R-type (ALU)
                id_is_rtype = 1; id_reg_we = 1; 
                // Decode R-type ALU operation based on funct3 and funct7
                case ({id_funct7, id_funct3})
                    10'b0000000_000: id_alu_op = ALU_ADD;  // ADD
                    10'b0100000_000: id_alu_op = ALU_SUB;  // SUB
                    10'b0000000_001: id_alu_op = ALU_SLL;  // SLL(Shift Left Logical)
                    10'b0000000_010: id_alu_op = ALU_SLT;  // SLT(Set less than)
                    10'b0000000_011: id_alu_op = ALU_SLTU; // SLTU(Set less than unsigned)
                    10'b0000000_100: id_alu_op = ALU_XOR;  // XOR
                    10'b0000000_101: id_alu_op = ALU_SRL;  // SRL(Shift right logical)
                    10'b0100000_101: id_alu_op = ALU_SRA;  // SRA(Shift right arithemetic)
                    10'b0000000_110: id_alu_op = ALU_OR;   // OR
                    10'b0000000_111: id_alu_op = ALU_AND;  // AND
                    default: id_alu_op = ALU_ADD;
                endcase
            end
            7'b0010011: begin // I-type ALU
                id_is_itype_alu = 1; id_reg_we = 1; 
                // Decode I-type ALU operation based on funct3 (shift instructions check funct7)
                case (id_funct3)
                    3'b000: id_alu_op = ALU_ADD;  // ADDI
                    3'b001: id_alu_op = ALU_SLL;  // SLLI
                    3'b010: id_alu_op = ALU_SLT;  // SLTI
                    3'b011: id_alu_op = ALU_SLTU; // SLTIU
                    3'b100: id_alu_op = ALU_XOR;  // XORI
                    3'b101: begin 
                        if (id_funct7[5] == 1'b0) id_alu_op = ALU_SRL; // SRLI
                        else id_alu_op = ALU_SRA; // SRAI
                    end
                    3'b110: id_alu_op = ALU_OR;   // ORI
                    3'b111: id_alu_op = ALU_AND;  // ANDI
                    default: id_alu_op = ALU_ADD;
                endcase
            end
            7'b0000011: begin id_is_load = 1; id_reg_we = 1; id_alu_op = ALU_ADD; end // Load
            7'b0100011: begin id_is_store = 1; id_alu_op = ALU_ADD; end // Store
            7'b1100011: id_is_branch = 1; // Branch
            7'b1101111: begin id_is_jal = 1; id_reg_we = 1; id_alu_op = ALU_ADD; end // JAL
            7'b1100111: begin id_is_jalr = 1; id_reg_we = 1; id_alu_op = ALU_ADD; end // JALR
            7'b0110111: begin id_reg_we = 1; id_alu_op = ALU_ADD; end // LUI
            7'b0010111: begin id_reg_we = 1; id_alu_op = ALU_ADD; end // AUIPC
            default: ;
        endcase
    end
    
    // -----------------------------------------------------------------
    //  HAZARD DETECTION UNIT (ID Stage)
    // -----------------------------------------------------------------
    always_comb begin
        // Default, No stall, no bubble
        pc_stall = 1'b0;
        id_ex_bubble = 1'b0;
        
        /* Load-Use Hazard Detection: 
        If the instruction in EX is a LOAD (id_ex_is_load)
         AND the Load's destination register (id_ex_rd) is needed by the ID instruction (id_rs1 or id_rs2)
        */
        if (id_ex_is_load && (id_ex_rd != 5'b0)) begin
            if ( (id_rs1 == id_ex_rd) || 
                (id_rs2 == id_ex_rd && (id_is_rtype || id_is_store || id_is_branch) ) )
            begin
                pc_stall = 1'b1;      // Freeze PC and IF/ID
                id_ex_bubble = 1'b1; // Insert NOP/Bubble into ID/EX
            end
        end
    end


    // -----------------------------------------------------------------
    //  FORWARDING UNIT 
    // -----------------------------------------------------------------
    
    always_comb begin
        forward_a = 2'b00; 
        forward_b = 2'b00;

        // --- Forwarding A (for RS1) ---
        // 1. EX/MEM -> EX Forwarding (Newest)
        if (ex_mem_reg_we && (ex_mem_rd != 5'b0) && (id_ex_rs1 == ex_mem_rd)) begin
            forward_a = 2'b01; 
        end
        // 2. MEM/WB -> EX Forwarding (Older, only if EX/MEM doesn't match)
        else if (mem_wb_reg_we && (mem_wb_rd != 5'b0) && (id_ex_rs1 == mem_wb_rd)) begin
            forward_a = 2'b10; 
        end
        
        // --- Forwarding B (for RS2) ---
        // 3. EX/MEM -> EX Forwarding (Newest)
        if (ex_mem_reg_we && (ex_mem_rd != 5'b0) && (id_ex_rs2 == ex_mem_rd)) begin
            forward_b = 2'b01; 
        end
        // 4. MEM/WB -> EX Forwarding (Older, only if EX/MEM doesn't match)
        else if (mem_wb_reg_we && (mem_wb_rd != 5'b0) && (id_ex_rs2 == mem_wb_rd)) begin
            forward_b = 2'b10; 
        end
    end
    
    // ID/EX Register Update (Includes NOP Insertion for Stall)
    always_ff @(posedge clk or posedge rst_p) begin
        if (rst_p) begin
            id_ex_instr    <= 32'b0;
            id_ex_pc       <= 32'b0;
            id_ex_rdata1   <= 32'b0;
            id_ex_rdata2   <= 32'b0;
            id_ex_imm      <= 32'b0;
            id_ex_alu_op   <= ALU_ADD;
            id_ex_reg_we   <= 1'b0;
            id_ex_is_load  <= 1'b0;
            id_ex_is_store <= 1'b0;
            id_ex_is_branch <= 1'b0;
            id_ex_is_jal   <= 1'b0;
            id_ex_is_jalr  <= 1'b0;
            id_ex_is_rtype <= 1'b0;
            id_ex_is_itype_alu <= 1'b0;
            id_ex_rs1      <= 5'b0; 
            id_ex_rs2      <= 5'b0;
            id_ex_rd       <= 5'b0;
        end else if (id_ex_bubble) begin // If hazard detected, insert NOP
            id_ex_instr    <= 32'b0;
            id_ex_reg_we   <= 1'b0; // Forces NOP
            id_ex_is_load  <= 1'b0; 
            id_ex_is_store <= 1'b0;
            id_ex_is_branch <= 1'b0;
            id_ex_is_jal   <= 1'b0;
            id_ex_is_jalr  <= 1'b0;
            id_ex_alu_op   <= ALU_ADD;
            id_ex_pc       <= 32'b0;
            id_ex_rd       <= 5'b0;
            // Other fields don't matter as reg_we=0
        end else begin // Normal data transfer
            id_ex_instr    <= if_id_instr;
            id_ex_pc       <= if_id_pc;
            id_ex_rdata1   <= id_rdata1; 
            id_ex_rdata2   <= id_rdata2; 
            
            if (id_is_store) id_ex_imm <= id_imm_s;
            else if (id_is_branch) id_ex_imm <= id_imm_b;
            else if (id_is_jal) id_ex_imm <= id_imm_j;
            else if (id_opcode == 7'b0110111 || id_opcode == 7'b0010111) id_ex_imm <= id_imm_u_shifted;
            else id_ex_imm <= id_imm_i; // I-type, JALR uses I-type
            
            id_ex_alu_op   <= id_alu_op;
            id_ex_reg_we   <= id_reg_we;
            id_ex_is_load  <= id_is_load;
            id_ex_is_store <= id_is_store;
            id_ex_is_branch <= id_is_branch;
            id_ex_is_jal   <= id_is_jal;
            id_ex_is_jalr  <= id_is_jalr;
            id_ex_is_rtype <= id_is_rtype;
            id_ex_is_itype_alu <= id_is_itype_alu;
            id_ex_rs1      <= id_rs1; 
            id_ex_rs2      <= id_rs2;
            id_ex_rd       <= id_rd;
        end
    end


    // =========================================================================
    // STAGE 3: EXECUTE (EX)
    // =========================================================================
    
    
    logic [31:0] ex_fwd_data_mem_wb; 
    logic [31:0] ex_fwd_data_ex_mem; 

    // EX Stage Forwarding Data Sources
    assign ex_fwd_data_ex_mem = ex_mem_alu_out;
    
    assign ex_fwd_data_mem_wb = (mem_wb_is_load) ? mem_wb_mem_rdata :  
                                (mem_wb_is_jal)  ? mem_wb_pc_plus_4 :  
                                                   mem_wb_alu_out;
    
    // ALU Input Selection with Forwarding
    logic [31:0] ex_alu_a_fwd, ex_alu_b_fwd;
    //dmem out declaration
    assign dmem_addr = ex_mem_alu_out[31:2]; // word-address for data memory
    assign dmem_addr_ip = ex_mem_alu_out[11:2];
    always_comb begin
        case (forward_a)
            2'b01: ex_alu_a_fwd = ex_fwd_data_ex_mem; 
            2'b10: ex_alu_a_fwd = ex_fwd_data_mem_wb; 
            default: ex_alu_a_fwd = id_ex_rdata1;     
        endcase
    end
    
    always_comb begin
        case (forward_b)
            2'b01: ex_alu_b_fwd = ex_fwd_data_ex_mem;
            2'b10: ex_alu_b_fwd = ex_fwd_data_mem_wb;
            default: ex_alu_b_fwd = id_ex_rdata2;
        endcase
    end
    
    // ALU Input Selection
    logic [31:0] ex_alu_a, ex_alu_b;
    always_comb begin
        ex_alu_a = ex_alu_a_fwd; 
        ex_alu_b = ex_alu_b_fwd;

        // I/S/JALR-type instructions use immediate as second operand
        if (id_ex_is_itype_alu || id_ex_is_load || id_ex_is_store || id_ex_is_jalr) begin
            ex_alu_b = id_ex_imm;
        end 
        
        // Special case for AUIPC/LUI (PC+Immediate or 0+Immediate)
        if (id_ex_instr[6:0] == 7'b0010111) begin // AUIPC
            ex_alu_a = id_ex_pc;
            ex_alu_b = id_ex_imm;
        end else if (id_ex_instr[6:0] == 7'b0110111) begin // LUI
            ex_alu_a = 32'b0;
            ex_alu_b = id_ex_imm;
        end
    end
    
    // ALU Execution 
    logic [31:0] ex_alu_out;
    always_comb begin
        ex_alu_out = 32'hX; // Default 

        unique case (id_ex_alu_op)
            ALU_ADD:  ex_alu_out = ex_alu_a + ex_alu_b; //ADD
            ALU_SUB:  ex_alu_out = ex_alu_a - ex_alu_b; //SUBTRACT
            ALU_SLL:  ex_alu_out = ex_alu_a << ex_alu_b[4:0]; //SLL
            ALU_SLT:  ex_alu_out = ($signed(ex_alu_a) < $signed(ex_alu_b)) ? 32'd1 : 32'd0;//SLT 
            ALU_SLTU: ex_alu_out = (ex_alu_a < ex_alu_b) ? 32'd1 : 32'd0; //SLTU
            ALU_XOR:  ex_alu_out = ex_alu_a ^ ex_alu_b;//XOR
            ALU_SRL:  ex_alu_out = ex_alu_a >> ex_alu_b[4:0];//SRL
            ALU_SRA:  ex_alu_out = $signed(ex_alu_a) >>> ex_alu_b[4:0]; // SRA
            ALU_OR:   ex_alu_out = ex_alu_a | ex_alu_b;//OR(Bitwise)
            ALU_AND:  ex_alu_out = ex_alu_a & ex_alu_b;//AND(Bitwise)
            default: ex_alu_out = 32'hX;//NOP
        endcase
    end
    logic branch_condition_met;
    
    logic [2:0] funct3 = id_ex_instr[14:12];
    // -----------------------------------------------------------------
    //  CONTROL HAZARD RESOLUTION UNIT (EX Stage) 
    // -----------------------------------------------------------------
    always_comb begin
        ex_branch_taken = 1'b0;
        ex_branch_target = id_ex_pc + 4; // Default target
        branch_condition_met = 1'b0;
        // 1. Jumps (Always Taken)
        if (id_ex_is_jal) begin
            ex_branch_taken = 1'b1;
            // JAL target is PC + Immediate (which is id_ex_imm)
            ex_branch_target = id_ex_pc + id_ex_imm; 
        end 
        else if (id_ex_is_jalr) begin
            ex_branch_taken = 1'b1;
            // JALR target is (rs1 + Immediate) & ~1
            ex_branch_target = (ex_alu_a_fwd + id_ex_imm) & 32'hFFFFFFFE; 
        end
        
        // 2. Conditional Branches (Resolved based on ALU inputs)
        else if (id_ex_is_branch) begin

            unique case (funct3)
                3'b000: branch_condition_met = (ex_alu_a_fwd == ex_alu_b_fwd); // BEQ(Branch Equal)
                3'b001: branch_condition_met = (ex_alu_a_fwd != ex_alu_b_fwd); // BNE(Branch Not equal)
                3'b100: branch_condition_met = ($signed(ex_alu_a_fwd) < $signed(ex_alu_b_fwd)); // BLT(Branch Less than)
                3'b101: branch_condition_met = ($signed(ex_alu_a_fwd) >= $signed(ex_alu_b_fwd)); // BGE(Branch greater than or equal)
                3'b110: branch_condition_met = (ex_alu_a_fwd < ex_alu_b_fwd); // BLTU(Branch less than unsigned)
                3'b111: branch_condition_met = (ex_alu_a_fwd >= ex_alu_b_fwd); // BGEU(Branch greater than or equal unsigned)
                default: branch_condition_met = 1'b0;
            endcase
            
            if (branch_condition_met) begin
                ex_branch_taken = 1'b1;
                // Branch target is PC + Immediate (which is id_ex_imm)
                ex_branch_target = id_ex_pc + id_ex_imm; 
            end
        end
    end
 
    // EX/MEM Register Update
    always_ff @(posedge clk or posedge rst_p) begin
        if (rst_p) begin
            ex_mem_alu_out <= 32'b0;
            ex_mem_wdata   <= 32'b0;
            ex_mem_rd      <= 5'b0;
            ex_mem_reg_we  <= 1'b0;
            ex_mem_mem_we  <= 1'b0;
            ex_mem_is_load <= 1'b0;
            ex_mem_is_jal  <= 1'b0;
            ex_mem_pc_plus_4 <= 32'b0;
        end else begin
            ex_mem_alu_out <= ex_alu_out;
            
            // Data for store comes from RS2, using forwarded value
            ex_mem_wdata   <= ex_alu_b_fwd; 
            
            ex_mem_rd      <= id_ex_rd;

            ex_mem_reg_we  <= id_ex_reg_we;
            ex_mem_mem_we  <= id_ex_is_store; 
            ex_mem_is_load <= id_ex_is_load;
            ex_mem_is_jal  <= id_ex_is_jal | id_ex_is_jalr;
            ex_mem_pc_plus_4 <= id_ex_pc + 4;
        end
    end


    // =========================================================================
    // STAGE 4: MEMORY ACCESS (MEM)
    // =========================================================================
    
    // Data Memory Read 
    wire [31:0] mem_dmem_rdata =dmem_dout;

    // Data Memory Write (Synchronous)
    always_ff @(posedge clk) begin
        if (ex_mem_mem_we) begin
            dmem[$clog2(DMEM_WORDS)'(ex_mem_alu_out[31:2])] <= ex_mem_wdata;
        end
    end
    
    // MEM/WB Register Update
    always_ff @(posedge clk or posedge rst_p) begin
        if (rst_p) begin
            mem_wb_alu_out   <= 32'b0;
            mem_wb_mem_rdata <= 32'b0;
            mem_wb_pc_plus_4 <= 32'b0;
            mem_wb_rd        <= 5'b0;
            mem_wb_reg_we    <= 1'b0;
            mem_wb_is_load   <= 1'b0;
            mem_wb_is_jal    <= 1'b0;
        end else begin
            mem_wb_alu_out   <= ex_mem_alu_out;
            mem_wb_mem_rdata <= mem_dmem_rdata;
            mem_wb_pc_plus_4 <= ex_mem_pc_plus_4;
            mem_wb_rd        <= ex_mem_rd;
            mem_wb_reg_we    <= ex_mem_reg_we;
            mem_wb_is_load   <= ex_mem_is_load;
            mem_wb_is_jal    <= ex_mem_is_jal;
        end
    end

    // =========================================================================
    // STAGE 5: WRITE BACK (WB)
    // =========================================================================
    
    // WB Data Selection 
    wire [31:0] wb_data;
    assign wb_data = (mem_wb_is_load) ? mem_wb_mem_rdata :  
                     (mem_wb_is_jal)  ? mem_wb_pc_plus_4 :  
                                        mem_wb_alu_out;    

    // Register File Write (Synchronous)
    always_ff @(posedge clk) begin
        if (mem_wb_reg_we && (mem_wb_rd != 5'b0)) begin
            regs[mem_wb_rd] <= wb_data;
        end
        else regs[0] <= 32'b0;
    end
     
endmodule
